* SPICE3 file created from clr.ext - technology: scmos

.option scale=1u

M1000 a_33_50# a_n13_27# myVdd Vdd pfet w=7 l=3
+ ad=63 pd=32 as=228 ps=110 
M1001 myVdd myIn a_33_50# Vdd pfet w=7 l=3
+ ad=0 pd=0 as=0 ps=0 
M1002 myOut a_33_50# myVdd Vdd pfet w=7 l=3
+ ad=63 pd=32 as=0 ps=0 
M1003 a_n13_27# myClr myVdd Vdd pfet w=5 l=3
+ ad=55 pd=32 as=0 ps=0 
M1004 a_n13_27# myClr myGnd Gnd nfet w=4 l=3
+ ad=48 pd=32 as=152 ps=90 
M1005 a_33_8# a_n13_27# myGnd Gnd nfet w=6 l=3
+ ad=54 pd=30 as=0 ps=0 
M1006 a_33_50# myIn a_33_8# Gnd nfet w=6 l=3
+ ad=42 pd=26 as=0 ps=0 
M1007 myOut a_33_50# myGnd Gnd nfet w=6 l=3
+ ad=72 pd=36 as=0 ps=0 
C0 myGnd gnd! 24.7fF
C1 myOut gnd! 8.3fF
C2 myClr gnd! 10.3fF
C3 myVdd gnd! 24.2fF
C4 a_33_50# gnd! 25.2fF
C5 myIn gnd! 33.1fF
C6 a_n13_27# gnd! 23.5fF
