* SPICE3 file created from antistrofeas3.ext - technology: scmos

.option scale=1u

M1000 out1 Vout inverter_2/Vdd Vdd pfet w=6 l=2
+ ad=52 pd=44 as=26 ps=22 
M1001 out1 Vout GND Gnd nfet w=3 l=2
+ ad=38 pd=36 as=57 ps=54 
M1002 out1 Vout Vdd Vdd pfet w=6 l=2
+ ad=0 pd=0 as=52 ps=44 
M1003 out1 Vout GND Gnd nfet w=3 l=2
+ ad=0 pd=0 as=0 ps=0 
M1004 Vout Vin Vdd Vdd pfet w=6 l=2
+ ad=26 pd=22 as=0 ps=0 
M1005 Vout Vin GND Gnd nfet w=3 l=2
+ ad=19 pd=18 as=0 ps=0 
C0 Vin gnd! 5.2fF
C1 Vdd gnd! 17.6fF
C2 out1 gnd! 11.6fF
C3 Vout gnd! 25.8fF


.include ../usc-spice.usc-spice

Vgnd1 GND 0 DC 0V
Vgnd2 gnd! 0 DC 0V
VVdd Vdd 0 DC 2.8V
Vin Vin 0 pulse(0 2.8 0ns 0.1ns 0.1ns 10ns 20ns)
.tran 5ns 40ns
.probe
.control
run
plot Vin out1+4
.endc
.end