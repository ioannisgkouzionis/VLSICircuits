* SPICE3 file created from poly_delay12.ext - technology: scmos

M1000 output inverter_11/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=312p ps=264u 
M1001 output inverter_11/in.t1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=228p ps=216u 
M1002 inverter_11/in.t0 inverter_9/out.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1003 inverter_11/in.t0 inverter_9/out.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1004 inverter_9/out.t0 inverter_9/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1005 inverter_9/out.t0 inverter_9/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1006 inverter_9/in.t0 inverter_8/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1007 inverter_9/in.t0 inverter_8/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1008 inverter_8/in.t0 inverter_7/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1009 inverter_8/in.t0 inverter_7/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1010 inverter_7/in.t0 inverter_6/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1011 inverter_7/in.t0 inverter_6/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1012 inverter_6/in.t0 inverter_5/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1013 inverter_6/in.t0 inverter_5/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1014 inverter_5/in.t0 inverter_4/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1015 inverter_5/in.t0 inverter_4/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1016 inverter_4/in.t0 inverter_3/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1017 inverter_4/in.t0 inverter_3/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1018 inverter_3/in.t0 inverter_2/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1019 inverter_3/in.t0 inverter_2/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1020 inverter_2/in.t0 inverter_1/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1021 inverter_2/in.t0 inverter_1/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1022 inverter_1/in.t0 input Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1023 inverter_1/in.t0 input GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
R0 inverter_11/in.t0 inverter_11/in.t1 43400
R1 inverter_9/out.t0 inverter_9/out.t1 43388
R2 inverter_9/in.t0 inverter_9/in.t1 43400
R3 inverter_8/in.t0 inverter_8/in.t1 43388
R4 inverter_7/in.t0 inverter_7/in.t1 43400
R5 inverter_6/in.t0 inverter_6/in.t1 43388
R6 inverter_5/in.t0 inverter_5/in.t1 43400
R7 inverter_4/in.t0 inverter_4/in.t1 43388
R8 inverter_3/in.t0 inverter_3/in.t1 43400
R9 inverter_2/in.t0 inverter_2/in.t1 43388
R10 inverter_1/in.t0 inverter_1/in.t1 43400
C0 inverter_1/in.t1 gnd! 430.5fF
C1 inverter_1/in.t0 gnd! 442.2fF
C2 inverter_2/in.t1 gnd! 430.4fF
C3 inverter_2/in.t0 gnd! 442.1fF
C4 inverter_3/in.t1 gnd! 430.5fF
C5 inverter_3/in.t0 gnd! 442.2fF
C6 inverter_4/in.t1 gnd! 430.4fF
C7 inverter_4/in.t0 gnd! 442.1fF
C8 inverter_5/in.t1 gnd! 430.5fF
C9 inverter_5/in.t0 gnd! 442.2fF
C10 inverter_6/in.t1 gnd! 430.4fF
C11 inverter_6/in.t0 gnd! 442.1fF
C12 inverter_7/in.t1 gnd! 430.5fF
C13 inverter_7/in.t0 gnd! 442.2fF
C14 inverter_8/in.t1 gnd! 430.4fF
C15 inverter_8/in.t0 gnd! 442.1fF
C16 inverter_9/in.t1 gnd! 430.4fF
C17 inverter_9/in.t0 gnd! 442.1fF
C18 inverter_9/out.t1 gnd! 430.4fF
C19 inverter_9/out.t0 gnd! 442.1fF
C20 inverter_11/in.t1 gnd! 430.5fF
C21 inverter_11/in.t0 gnd! 442.2fF
C22 input gnd! 5.2fF
C23 Vdd gnd! 5658.1fF

.include ../usc-spice.usc-spice

Vgnd1 GND 0 DC 0VZ
Vgnd2 gnd! 0 DC 0V
VVdd Vdd 0 DC 2.8V
Vin input 0 pulse(0 2.8 0ns 0.1ns 0.1ns 5000ns 10000ns)
.tran 5ns 20000ns
.probe
.control
run
plot input output+4
.endc
.end

