magic
tech scmos
timestamp 1477223331
<< nwell >>
rect -26 -2 36 8
rect -33 -60 57 -50
<< polysilicon >>
rect -13 7 -9 19
rect 19 7 23 19
rect -13 -9 -9 1
rect 19 -9 23 1
rect -13 -32 -9 -15
rect 3 -32 7 -13
rect 19 -32 23 -15
rect 38 -32 42 -13
rect -13 -50 -9 -38
rect 3 -50 7 -38
rect 19 -50 23 -38
rect 38 -50 42 -38
rect -13 -65 -9 -57
rect 3 -65 7 -57
rect 19 -65 23 -57
rect 38 -65 42 -57
<< ndiffusion >>
rect -20 -10 -13 -9
rect -20 -14 -19 -10
rect -15 -14 -13 -10
rect -20 -15 -13 -14
rect -9 -10 -1 -9
rect -9 -14 -7 -10
rect -3 -14 -1 -10
rect -9 -15 -1 -14
rect 13 -10 19 -9
rect 13 -14 14 -10
rect 18 -14 19 -10
rect 13 -15 19 -14
rect 23 -10 31 -9
rect 23 -14 25 -10
rect 29 -14 31 -10
rect 23 -15 31 -14
rect -30 -33 -13 -32
rect -30 -37 -19 -33
rect -15 -37 -13 -33
rect -30 -38 -13 -37
rect -9 -33 3 -32
rect -9 -37 -5 -33
rect -1 -37 3 -33
rect -9 -38 3 -37
rect 7 -33 19 -32
rect 7 -37 11 -33
rect 15 -37 19 -33
rect 7 -38 19 -37
rect 23 -33 38 -32
rect 23 -37 29 -33
rect 33 -37 38 -33
rect 23 -38 38 -37
rect 42 -33 54 -32
rect 42 -37 49 -33
rect 53 -37 54 -33
rect 42 -38 54 -37
<< pdiffusion >>
rect -20 6 -13 7
rect -20 2 -19 6
rect -15 2 -13 6
rect -20 1 -13 2
rect -9 6 -2 7
rect -9 2 -7 6
rect -3 2 -2 6
rect -9 1 -2 2
rect 12 6 19 7
rect 12 2 13 6
rect 17 2 19 6
rect 12 1 19 2
rect 23 6 30 7
rect 23 2 25 6
rect 29 2 30 6
rect 23 1 30 2
rect -32 -52 -13 -50
rect -32 -56 -19 -52
rect -15 -56 -13 -52
rect -32 -57 -13 -56
rect -9 -52 3 -50
rect -9 -56 -4 -52
rect 0 -56 3 -52
rect -9 -57 3 -56
rect 7 -57 19 -50
rect 23 -52 38 -50
rect 23 -56 29 -52
rect 33 -56 38 -52
rect 23 -57 38 -56
rect 42 -52 54 -50
rect 42 -56 49 -52
rect 53 -56 54 -52
rect 42 -57 54 -56
<< metal1 >>
rect -41 9 70 14
rect -19 6 -15 9
rect 13 6 17 9
rect -7 -3 -3 2
rect 25 -2 29 2
rect -7 -6 7 -3
rect -7 -10 -3 -6
rect 3 -9 7 -6
rect 25 -6 42 -2
rect 25 -10 29 -6
rect 38 -9 42 -6
rect -19 -17 -15 -14
rect 14 -17 18 -14
rect -35 -22 53 -17
rect -19 -33 -15 -22
rect -5 -30 33 -27
rect -5 -33 -1 -30
rect 29 -33 33 -30
rect 49 -33 53 -22
rect 11 -40 15 -37
rect -31 -43 15 -40
rect -31 -44 0 -43
rect -4 -52 0 -44
rect 66 -46 70 9
rect 29 -49 70 -46
rect 29 -52 33 -49
rect -19 -65 -15 -56
rect 49 -65 53 -56
rect -19 -68 53 -65
<< ntransistor >>
rect -13 -15 -9 -9
rect 19 -15 23 -9
rect -13 -38 -9 -32
rect 3 -38 7 -32
rect 19 -38 23 -32
rect 38 -38 42 -32
<< ptransistor >>
rect -13 1 -9 7
rect 19 1 23 7
rect -13 -57 -9 -50
rect 3 -57 7 -50
rect 19 -57 23 -50
rect 38 -57 42 -50
<< polycontact >>
rect 3 -13 7 -9
rect 38 -13 42 -9
<< ndcontact >>
rect -19 -14 -15 -10
rect -7 -14 -3 -10
rect 14 -14 18 -10
rect 25 -14 29 -10
rect -19 -37 -15 -33
rect -5 -37 -1 -33
rect 11 -37 15 -33
rect 29 -37 33 -33
rect 49 -37 53 -33
<< pdcontact >>
rect -19 2 -15 6
rect -7 2 -3 6
rect 13 2 17 6
rect 25 2 29 6
rect -19 -56 -15 -52
rect -4 -56 0 -52
rect 29 -56 33 -52
rect 49 -56 53 -52
<< labels >>
rlabel metal1 -36 11 -36 11 1 myVdd
rlabel polysilicon -11 17 -11 17 5 myIna
rlabel polysilicon 21 16 21 16 5 myInb
rlabel metal1 -30 -20 -30 -20 1 myGnd
rlabel metal1 -28 -42 -28 -42 1 myOut
<< end >>
