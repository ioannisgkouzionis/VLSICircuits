magic
tech scmos
timestamp 1477231015
<< nwell >>
rect -88 66 -26 76
rect 15 66 77 76
rect -109 0 -19 10
rect 8 0 98 10
<< polysilicon >>
rect -75 75 -71 87
rect -43 75 -39 87
rect 28 75 32 77
rect 60 75 64 87
rect -75 59 -71 69
rect -43 59 -39 69
rect 28 59 32 69
rect 60 59 64 69
rect -94 36 -90 55
rect -75 36 -71 53
rect -59 36 -55 55
rect -43 36 -39 53
rect 28 36 32 53
rect 44 36 48 55
rect 60 36 64 53
rect 79 36 83 55
rect -94 10 -90 30
rect -75 10 -71 30
rect -59 10 -55 30
rect -43 10 -39 30
rect 28 27 32 30
rect 28 10 32 22
rect 44 10 48 30
rect 60 10 64 30
rect 79 10 83 30
rect -94 -5 -90 3
rect -75 -5 -71 3
rect -59 -5 -55 3
rect -43 -5 -39 3
rect 28 -5 32 3
rect 44 -5 48 3
rect 60 -5 64 3
rect 79 -5 83 3
<< ndiffusion >>
rect -83 58 -75 59
rect -83 54 -81 58
rect -77 54 -75 58
rect -83 53 -75 54
rect -71 58 -65 59
rect -71 54 -70 58
rect -66 54 -65 58
rect -71 53 -65 54
rect -51 58 -43 59
rect -51 54 -49 58
rect -45 54 -43 58
rect -51 53 -43 54
rect -39 58 -32 59
rect -39 54 -37 58
rect -33 54 -32 58
rect -39 53 -32 54
rect 21 58 28 59
rect 21 54 22 58
rect 26 54 28 58
rect 21 53 28 54
rect 32 58 40 59
rect 32 54 34 58
rect 38 54 40 58
rect 32 53 40 54
rect 54 58 60 59
rect 54 54 55 58
rect 59 54 60 58
rect 54 53 60 54
rect 64 58 72 59
rect 64 54 66 58
rect 70 54 72 58
rect 64 53 72 54
rect -106 35 -94 36
rect -106 31 -105 35
rect -101 31 -94 35
rect -106 30 -94 31
rect -90 35 -75 36
rect -90 31 -85 35
rect -81 31 -75 35
rect -90 30 -75 31
rect -71 35 -59 36
rect -71 31 -67 35
rect -63 31 -59 35
rect -71 30 -59 31
rect -55 35 -43 36
rect -55 31 -51 35
rect -47 31 -43 35
rect -55 30 -43 31
rect -39 35 -22 36
rect -39 31 -37 35
rect -33 31 -22 35
rect -39 30 -22 31
rect 11 35 28 36
rect 11 31 22 35
rect 26 31 28 35
rect 11 30 28 31
rect 32 35 44 36
rect 32 31 36 35
rect 40 31 44 35
rect 32 30 44 31
rect 48 35 60 36
rect 48 31 52 35
rect 56 31 60 35
rect 48 30 60 31
rect 64 35 79 36
rect 64 31 70 35
rect 74 31 79 35
rect 64 30 79 31
rect 83 35 95 36
rect 83 31 90 35
rect 94 31 95 35
rect 83 30 95 31
<< pdiffusion >>
rect -82 74 -75 75
rect -82 70 -81 74
rect -77 70 -75 74
rect -82 69 -75 70
rect -71 74 -64 75
rect -71 70 -69 74
rect -65 70 -64 74
rect -71 69 -64 70
rect -50 74 -43 75
rect -50 70 -49 74
rect -45 70 -43 74
rect -50 69 -43 70
rect -39 74 -32 75
rect -39 70 -37 74
rect -33 70 -32 74
rect -39 69 -32 70
rect 21 74 28 75
rect 21 70 22 74
rect 26 70 28 74
rect 21 69 28 70
rect 32 74 39 75
rect 32 70 34 74
rect 38 70 39 74
rect 32 69 39 70
rect 53 74 60 75
rect 53 70 54 74
rect 58 70 60 74
rect 53 69 60 70
rect 64 74 71 75
rect 64 70 66 74
rect 70 70 71 74
rect 64 69 71 70
rect -106 8 -94 10
rect -106 4 -105 8
rect -101 4 -94 8
rect -106 3 -94 4
rect -90 8 -75 10
rect -90 4 -85 8
rect -81 4 -75 8
rect -90 3 -75 4
rect -71 3 -59 10
rect -55 8 -43 10
rect -55 4 -52 8
rect -48 4 -43 8
rect -55 3 -43 4
rect -39 8 -20 10
rect -39 4 -37 8
rect -33 4 -20 8
rect -39 3 -20 4
rect 9 8 28 10
rect 9 4 22 8
rect 26 4 28 8
rect 9 3 28 4
rect 32 8 44 10
rect 32 4 37 8
rect 41 4 44 8
rect 32 3 44 4
rect 48 3 60 10
rect 64 8 79 10
rect 64 4 70 8
rect 74 4 79 8
rect 64 3 79 4
rect 83 8 95 10
rect 83 4 90 8
rect 94 4 95 8
rect 83 3 95 4
<< metal1 >>
rect -122 77 111 82
rect -122 14 -118 77
rect -69 74 -65 77
rect -37 74 -33 77
rect 22 74 26 77
rect 54 74 58 77
rect -81 66 -77 70
rect -94 62 -77 66
rect -49 65 -45 70
rect -94 59 -90 62
rect -81 58 -77 62
rect -59 62 -45 65
rect -59 59 -55 62
rect -49 58 -45 62
rect 34 65 38 70
rect 66 66 70 70
rect 34 62 48 65
rect 34 58 38 62
rect -70 51 -66 54
rect -37 51 -33 54
rect 44 59 48 62
rect 66 62 83 66
rect 66 58 70 62
rect 79 59 83 62
rect 22 51 26 54
rect 55 51 59 54
rect -105 46 94 51
rect -105 35 -101 46
rect -85 38 -47 41
rect -85 35 -81 38
rect -51 35 -47 38
rect -37 35 -33 46
rect 22 35 26 46
rect 36 38 74 41
rect 36 35 40 38
rect 70 35 74 38
rect 90 35 94 46
rect -67 27 -63 31
rect -67 22 28 27
rect -122 11 -81 14
rect -85 8 -81 11
rect -52 8 -48 22
rect 52 14 56 31
rect 107 14 111 77
rect 1 11 56 14
rect 70 11 111 14
rect -105 -5 -101 4
rect -37 -5 -33 4
rect -105 -8 -33 -5
rect 1 -13 5 11
rect 37 8 41 11
rect 70 8 74 11
rect 22 -5 26 4
rect 90 -5 94 4
rect 22 -8 94 -5
<< ntransistor >>
rect -75 53 -71 59
rect -43 53 -39 59
rect 28 53 32 59
rect 60 53 64 59
rect -94 30 -90 36
rect -75 30 -71 36
rect -59 30 -55 36
rect -43 30 -39 36
rect 28 30 32 36
rect 44 30 48 36
rect 60 30 64 36
rect 79 30 83 36
<< ptransistor >>
rect -75 69 -71 75
rect -43 69 -39 75
rect 28 69 32 75
rect 60 69 64 75
rect -94 3 -90 10
rect -75 3 -71 10
rect -59 3 -55 10
rect -43 3 -39 10
rect 28 3 32 10
rect 44 3 48 10
rect 60 3 64 10
rect 79 3 83 10
<< polycontact >>
rect -94 55 -90 59
rect -59 55 -55 59
rect 44 55 48 59
rect 79 55 83 59
rect 28 22 32 27
<< ndcontact >>
rect -81 54 -77 58
rect -70 54 -66 58
rect -49 54 -45 58
rect -37 54 -33 58
rect 22 54 26 58
rect 34 54 38 58
rect 55 54 59 58
rect 66 54 70 58
rect -105 31 -101 35
rect -85 31 -81 35
rect -67 31 -63 35
rect -51 31 -47 35
rect -37 31 -33 35
rect 22 31 26 35
rect 36 31 40 35
rect 52 31 56 35
rect 70 31 74 35
rect 90 31 94 35
<< pdcontact >>
rect -81 70 -77 74
rect -69 70 -65 74
rect -49 70 -45 74
rect -37 70 -33 74
rect 22 70 26 74
rect 34 70 38 74
rect 54 70 58 74
rect 66 70 70 74
rect -105 4 -101 8
rect -85 4 -81 8
rect -52 4 -48 8
rect -37 4 -33 8
rect 22 4 26 8
rect 37 4 41 8
rect 70 4 74 8
rect 90 4 94 8
<< labels >>
rlabel metal1 -115 79 -115 79 1 myVdd
rlabel metal1 -102 48 -102 48 1 myGnd
rlabel polysilicon -73 84 -73 84 5 myB
rlabel polysilicon -41 84 -41 84 5 myA
rlabel polysilicon 62 84 62 84 5 myCin
rlabel metal1 3 -7 3 -7 1 myOut
<< end >>
