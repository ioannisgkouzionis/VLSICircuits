magic
tech scmos
timestamp 1477235084
<< polysilicon >>
rect -13 32 3 34
rect 8 32 45 34
rect -13 31 45 32
rect -13 22 -10 31
rect 2 22 5 24
rect 20 22 24 24
rect 42 22 45 31
rect 51 22 55 32
rect 93 22 97 26
rect -13 -2 -10 15
rect 2 -2 5 15
rect 20 -2 24 15
rect 42 -2 45 15
rect 51 -2 55 15
rect 93 9 97 15
rect 95 3 97 9
rect 93 -1 97 3
rect -13 -12 -10 -9
rect 2 -14 5 -9
rect 20 -12 24 -9
rect 42 -12 45 -9
rect 51 -14 55 -9
rect 93 -12 97 -8
rect 2 -16 55 -14
<< ndiffusion >>
rect 83 -2 93 -1
rect -23 -3 -13 -2
rect -23 -8 -21 -3
rect -16 -8 -13 -3
rect -23 -9 -13 -8
rect -10 -3 2 -2
rect -10 -8 -6 -3
rect -1 -8 2 -3
rect -10 -9 2 -8
rect 5 -3 20 -2
rect 5 -8 9 -3
rect 14 -8 20 -3
rect 5 -9 20 -8
rect 24 -3 42 -2
rect 24 -8 31 -3
rect 36 -8 42 -3
rect 24 -9 42 -8
rect 45 -9 51 -2
rect 55 -3 68 -2
rect 55 -8 59 -3
rect 64 -8 68 -3
rect 83 -7 85 -2
rect 90 -7 93 -2
rect 83 -8 93 -7
rect 97 -2 108 -1
rect 97 -7 101 -2
rect 106 -7 108 -2
rect 97 -8 108 -7
rect 55 -9 68 -8
<< pdiffusion >>
rect -23 21 -13 22
rect -23 16 -21 21
rect -16 16 -13 21
rect -23 15 -13 16
rect -10 21 2 22
rect -10 16 -7 21
rect -2 16 2 21
rect -10 15 2 16
rect 5 21 20 22
rect 5 16 9 21
rect 14 16 20 21
rect 5 15 20 16
rect 24 21 42 22
rect 24 16 30 21
rect 35 16 42 21
rect 24 15 42 16
rect 45 15 51 22
rect 55 21 67 22
rect 55 16 59 21
rect 64 16 67 21
rect 55 15 67 16
rect 83 21 93 22
rect 83 16 85 21
rect 90 16 93 21
rect 83 15 93 16
rect 97 21 108 22
rect 97 16 101 21
rect 106 16 108 21
rect 97 15 108 16
<< metal1 >>
rect 21 44 44 49
rect 3 36 8 39
rect 20 28 24 39
rect -21 24 14 27
rect 30 27 35 44
rect 51 36 55 40
rect 30 24 90 27
rect -21 21 -16 24
rect 9 21 14 24
rect 30 21 35 24
rect 85 21 90 24
rect -7 13 -2 16
rect 59 13 64 16
rect -7 10 64 13
rect 59 9 64 10
rect 101 10 106 16
rect 59 3 91 9
rect 101 5 117 10
rect -6 0 64 3
rect -6 -3 -1 0
rect 59 -3 64 0
rect 101 -2 106 5
rect -21 -18 -16 -8
rect 9 -18 14 -8
rect -21 -21 14 -18
rect 31 -18 36 -8
rect 85 -18 90 -7
rect 31 -23 90 -18
rect 58 -27 66 -23
rect 49 -34 76 -27
<< ntransistor >>
rect -13 -9 -10 -2
rect 2 -9 5 -2
rect 20 -9 24 -2
rect 42 -9 45 -2
rect 51 -9 55 -2
rect 93 -8 97 -1
<< ptransistor >>
rect -13 15 -10 22
rect 2 15 5 22
rect 20 15 24 22
rect 42 15 45 22
rect 51 15 55 22
rect 93 15 97 22
<< polycontact >>
rect 3 32 8 36
rect 20 24 24 28
rect 51 32 55 36
rect 91 3 95 9
<< ndcontact >>
rect -21 -8 -16 -3
rect -6 -8 -1 -3
rect 9 -8 14 -3
rect 31 -8 36 -3
rect 59 -8 64 -3
rect 85 -7 90 -2
rect 101 -7 106 -2
<< pdcontact >>
rect -21 16 -16 21
rect -7 16 -2 21
rect 9 16 14 21
rect 30 16 35 21
rect 59 16 64 21
rect 85 16 90 21
rect 101 16 106 21
<< labels >>
rlabel metal1 33 46 33 46 5 myVdd
rlabel metal1 6 37 6 37 1 myB
rlabel metal1 22 37 22 37 1 myA
rlabel metal1 53 38 53 38 1 myCin
rlabel metal1 63 -30 63 -30 1 myGnd
rlabel metal1 113 7 113 7 7 myOut
<< end >>
