magic
tech scmos
timestamp 1415315269
<< polysilicon >>
rect 113 412 158 414
rect 112 380 126 382
rect 254 380 266 382
rect 196 355 201 357
rect 56 353 64 355
rect 69 313 90 315
rect -1 308 8 310
rect 133 310 135 315
rect 209 313 230 315
rect 133 308 148 310
rect 157 114 161 116
rect 32 111 34 114
rect 157 109 159 114
<< metal1 >>
rect 3 424 6 430
rect 75 427 146 430
rect 19 424 22 427
rect 75 415 78 427
rect 143 421 146 427
rect 202 414 205 426
rect 215 427 259 430
rect 215 415 218 427
rect 127 362 130 380
rect 267 360 270 378
rect 61 346 64 349
rect 199 348 202 351
rect 201 344 202 348
rect 12 308 15 311
rect 66 310 69 313
rect 152 307 155 310
rect 206 310 209 313
rect 32 102 35 107
rect 156 102 159 105
rect -3 9 32 12
rect 36 9 156 12
rect 160 9 268 12
<< metal2 >>
rect 23 427 201 430
rect 2 417 62 420
rect 127 347 130 358
rect 1 342 60 345
rect 127 344 197 347
rect 1 333 50 336
rect 121 333 190 336
rect 261 333 273 336
rect 1 324 23 327
rect 27 324 163 327
rect 167 324 273 327
rect 19 307 65 310
rect 159 307 205 310
rect 32 13 35 98
rect 156 13 159 98
<< polycontact >>
rect 126 380 130 384
rect 266 378 270 382
rect 60 349 64 353
rect 199 351 203 355
rect 65 313 69 317
rect 8 307 12 311
rect 205 313 209 317
rect 148 307 152 311
rect 31 107 35 111
rect 155 105 159 109
<< m2contact >>
rect 19 427 23 431
rect 62 416 66 420
rect 201 426 205 430
rect 127 358 131 362
rect 267 356 271 360
rect 60 342 64 346
rect 197 344 201 348
rect 50 333 54 337
rect 117 333 121 337
rect 190 332 194 336
rect 257 333 261 337
rect 23 323 27 327
rect 163 323 167 327
rect 15 307 19 311
rect 65 306 69 310
rect 155 307 159 311
rect 205 306 209 310
rect 31 98 35 102
rect 155 98 159 102
rect 32 9 36 13
rect 156 9 160 13
use shiftregistermodule  shiftregistermodule_0
timestamp 1415310808
transform 0 1 0 -1 0 316
box -108 0 296 133
use shiftregistermodule  shiftregistermodule_1
timestamp 1415310808
transform 0 1 140 -1 0 316
box -108 0 296 133
<< end >>
