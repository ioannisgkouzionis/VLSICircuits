* SPICE3 file created from poly_delay14.ext - technology: scmos

M1000 output inverter_13/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=26p pd=22u as=364p ps=308u 
M1001 output inverter_13/in.t1 GND Gnd nfet w=3u l=2u
+ ad=19p pd=18u as=266p ps=252u 
M1002 inverter_13/in.t0 inverter_12/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1003 inverter_13/in.t0 inverter_12/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1004 inverter_12/in.t0 inverter_11/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1005 inverter_12/in.t0 inverter_11/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1006 inverter_11/in.t0 inverter_9/out.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1007 inverter_11/in.t0 inverter_9/out.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1008 inverter_9/out.t0 inverter_9/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1009 inverter_9/out.t0 inverter_9/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1010 inverter_9/in.t0 inverter_8/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1011 inverter_9/in.t0 inverter_8/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1012 inverter_8/in.t0 inverter_7/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1013 inverter_8/in.t0 inverter_7/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1014 inverter_7/in.t0 inverter_6/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1015 inverter_7/in.t0 inverter_6/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1016 inverter_6/in.t0 inverter_5/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1017 inverter_6/in.t0 inverter_5/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1018 inverter_5/in.t0 inverter_4/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1019 inverter_5/in.t0 inverter_4/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1020 inverter_4/in.t0 inverter_3/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1021 inverter_4/in.t0 inverter_3/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1022 inverter_3/in.t0 inverter_2/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1023 inverter_3/in.t0 inverter_2/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1024 inverter_2/in.t0 inverter_1/in.t1 Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1025 inverter_2/in.t0 inverter_1/in.t1 GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1026 inverter_1/in.t0 input Vdd Vdd pfet w=6u l=2u
+ ad=0p pd=0u as=0p ps=0u 
M1027 inverter_1/in.t0 input GND Gnd nfet w=3u l=2u
+ ad=0p pd=0u as=0p ps=0u 
R0 inverter_13/in.t0 inverter_13/in.t1 36671
R1 inverter_12/in.t0 inverter_12/in.t1 36755
R2 inverter_11/in.t0 inverter_11/in.t1 36671
R3 inverter_9/out.t0 inverter_9/out.t1 36731
R4 inverter_9/in.t0 inverter_9/in.t1 36707
R5 inverter_8/in.t0 inverter_8/in.t1 36707
R6 inverter_7/in.t0 inverter_7/in.t1 36707
R7 inverter_6/in.t0 inverter_6/in.t1 36707
R8 inverter_5/in.t0 inverter_5/in.t1 36707
R9 inverter_4/in.t0 inverter_4/in.t1 36707
R10 inverter_3/in.t0 inverter_3/in.t1 36707
R11 inverter_2/in.t0 inverter_2/in.t1 36707
R12 inverter_1/in.t0 inverter_1/in.t1 36707
C0 inverter_1/in.t1 gnd! 363.7fF
C1 inverter_1/in.t0 gnd! 375.5fF
C2 inverter_2/in.t1 gnd! 363.7fF
C3 inverter_2/in.t0 gnd! 375.5fF
C4 inverter_3/in.t1 gnd! 363.7fF
C5 inverter_3/in.t0 gnd! 375.5fF
C6 inverter_4/in.t1 gnd! 363.7fF
C7 inverter_4/in.t0 gnd! 375.5fF
C8 inverter_5/in.t1 gnd! 363.7fF
C9 inverter_5/in.t0 gnd! 375.5fF
C10 inverter_6/in.t1 gnd! 363.7fF
C11 inverter_6/in.t0 gnd! 375.5fF
C12 inverter_7/in.t1 gnd! 363.7fF
C13 inverter_7/in.t0 gnd! 375.5fF
C14 inverter_8/in.t1 gnd! 363.7fF
C15 inverter_8/in.t0 gnd! 375.5fF
C16 inverter_9/in.t1 gnd! 363.7fF
C17 inverter_9/in.t0 gnd! 375.5fF
C18 inverter_9/out.t1 gnd! 364.0fF
C19 inverter_9/out.t0 gnd! 375.7fF
C20 inverter_11/in.t1 gnd! 363.4fF
C21 inverter_11/in.t0 gnd! 375.1fF
C22 inverter_12/in.t1 gnd! 364.2fF
C23 inverter_12/in.t0 gnd! 375.9fF
C24 inverter_13/in.t1 gnd! 363.4fF
C25 inverter_13/in.t0 gnd! 375.1fF
C26 input gnd! 6.2fF
C27 Vdd gnd! 5659.0fF

.include ../usc-spice.usc-spice

Vgnd1 GND 0 DC 0VZ
Vgnd2 gnd! 0 DC 0V
VVdd Vdd 0 DC 2.8V
Vin input 0 pulse(0 2.8 0ns 0.1ns 0.1ns 5000ns 10000ns)
.tran 5ns 20000ns
.probe
.control
run
plot input output+4
.endc
.end
