* SPICE3 file created from dff2.ext - technology: scmos

.option scale=1u

M1000 not_0/myA myClk myVdd Vdd pfet w=5 l=3
+ ad=55 pd=32 as=1008 ps=552 
M1001 not_0/myA myClk myGnd Gnd nfet w=4 l=3
+ ad=48 pd=32 as=724 ps=480 
M1002 not_0/myOut not_0/myA myVdd Vdd pfet w=5 l=3
+ ad=55 pd=32 as=0 ps=0 
M1003 not_0/myOut not_0/myA myGnd Gnd nfet w=4 l=3
+ ad=48 pd=32 as=0 ps=0 
M1004 dff1_0/not_0/myA not_0/myOut myVdd Vdd pfet w=5 l=3
+ ad=55 pd=32 as=0 ps=0 
M1005 dff1_0/not_0/myA not_0/myOut myGnd Gnd nfet w=4 l=3
+ ad=48 pd=32 as=0 ps=0 
M1006 dff1_0/not_4/myOut dff1_0/not_0/myA myVdd Vdd pfet w=5 l=3
+ ad=55 pd=32 as=0 ps=0 
M1007 dff1_0/not_4/myOut dff1_0/not_0/myA myGnd Gnd nfet w=4 l=3
+ ad=48 pd=32 as=0 ps=0 
M1008 dff1_0/gate_0/myC dff1_0/not_0/myA myVdd Vdd pfet w=5 l=3
+ ad=55 pd=32 as=0 ps=0 
M1009 dff1_0/gate_0/myC dff1_0/not_0/myA myGnd Gnd nfet w=4 l=3
+ ad=48 pd=32 as=0 ps=0 
M1010 dff1_0/gate_1/myD dff1_0/not_2/myA myVdd Vdd pfet w=5 l=3
+ ad=110 pd=64 as=0 ps=0 
M1011 dff1_0/gate_1/myD dff1_0/not_2/myA myGnd Gnd nfet w=4 l=3
+ ad=96 pd=64 as=0 ps=0 
M1012 dff1_0/not_2/myA dff1_0/not_1/myA myVdd Vdd pfet w=5 l=3
+ ad=110 pd=64 as=0 ps=0 
M1013 dff1_0/not_2/myA dff1_0/not_1/myA myGnd Gnd nfet w=4 l=3
+ ad=96 pd=64 as=0 ps=0 
M1014 dff1_0/not_1/myA dff1_0/gate_1/a_3_46# dff1_0/gate_1/myD Vdd pfet w=5 l=3
+ ad=120 pd=68 as=0 ps=0 
M1015 dff1_0/not_1/myA dff1_0/not_0/myA dff1_0/gate_1/myD Gnd nfet w=4 l=3
+ ad=104 pd=68 as=0 ps=0 
M1016 dff1_0/gate_1/a_3_46# dff1_0/not_0/myA myVdd Vdd pfet w=5 l=3
+ ad=55 pd=32 as=0 ps=0 
M1017 dff1_0/gate_1/a_3_46# dff1_0/not_0/myA myGnd Gnd nfet w=4 l=3
+ ad=48 pd=32 as=0 ps=0 
M1018 dff1_0/not_1/myA dff1_0/gate_0/a_3_46# dff1_0/gate_0/myD Vdd pfet w=5 l=3
+ ad=0 pd=0 as=118 ps=64 
M1019 dff1_0/not_1/myA dff1_0/gate_0/myC dff1_0/gate_0/myD Gnd nfet w=4 l=3
+ ad=0 pd=0 as=120 ps=68 
M1020 dff1_0/gate_0/a_3_46# dff1_0/gate_0/myC myVdd Vdd pfet w=5 l=3
+ ad=55 pd=32 as=0 ps=0 
M1021 dff1_0/gate_0/a_3_46# dff1_0/gate_0/myC myGnd Gnd nfet w=4 l=3
+ ad=48 pd=32 as=0 ps=0 
M1022 dff1_0/clr_0/a_33_50# dff1_0/clr_0/a_n13_27# myVdd Vdd pfet w=7 l=3
+ ad=63 pd=32 as=0 ps=0 
M1023 myVdd myD dff1_0/clr_0/a_33_50# Vdd pfet w=7 l=3
+ ad=0 pd=0 as=0 ps=0 
M1024 dff1_0/gate_0/myD dff1_0/clr_0/a_33_50# myVdd Vdd pfet w=7 l=3
+ ad=0 pd=0 as=0 ps=0 
M1025 dff1_0/clr_0/a_n13_27# myClr myVdd Vdd pfet w=5 l=3
+ ad=55 pd=32 as=0 ps=0 
M1026 dff1_0/clr_0/a_n13_27# myClr myGnd Gnd nfet w=4 l=3
+ ad=48 pd=32 as=0 ps=0 
M1027 dff1_0/clr_0/a_33_8# dff1_0/clr_0/a_n13_27# myGnd Gnd nfet w=6 l=3
+ ad=54 pd=30 as=0 ps=0 
M1028 dff1_0/clr_0/a_33_50# myD dff1_0/clr_0/a_33_8# Gnd nfet w=6 l=3
+ ad=42 pd=26 as=0 ps=0 
M1029 dff1_0/gate_0/myD dff1_0/clr_0/a_33_50# myGnd Gnd nfet w=6 l=3
+ ad=0 pd=0 as=0 ps=0 
M1030 myOut1 dff1_0/a_n133_170# dff1_0/not_2/myA Vdd pfet w=5 l=3
+ ad=120 pd=68 as=0 ps=0 
M1031 myOut1 dff1_0/not_0/myA dff1_0/not_2/myA Gnd nfet w=4 l=3
+ ad=104 pd=68 as=0 ps=0 
M1032 dff1_0/a_n56_158# dff1_0/a_n81_156# myOut1 Vdd pfet w=5 l=3
+ ad=110 pd=64 as=0 ps=0 
M1033 myOut2 myOut1 myVdd Vdd pfet w=5 l=3
+ ad=55 pd=32 as=0 ps=0 
M1034 dff1_0/a_n56_158# dff1_0/not_4/myOut myOut1 Gnd nfet w=4 l=3
+ ad=96 pd=64 as=0 ps=0 
M1035 myOut2 myOut1 myGnd Gnd nfet w=4 l=3
+ ad=48 pd=32 as=0 ps=0 
M1036 dff1_0/a_n133_170# dff1_0/not_0/myA myVdd Vdd pfet w=5 l=3
+ ad=55 pd=32 as=0 ps=0 
M1037 myVdd dff1_0/not_4/myOut dff1_0/a_n81_156# Vdd pfet w=5 l=3
+ ad=0 pd=0 as=55 ps=32 
M1038 myVdd myOut2 dff1_0/a_n56_158# Vdd pfet w=5 l=3
+ ad=0 pd=0 as=0 ps=0 
M1039 dff1_0/a_n133_170# dff1_0/not_0/myA myGnd Gnd nfet w=4 l=3
+ ad=48 pd=32 as=0 ps=0 
M1040 myGnd dff1_0/not_4/myOut dff1_0/a_n81_156# Gnd nfet w=4 l=3
+ ad=0 pd=0 as=48 ps=32 
M1041 myGnd myOut2 dff1_0/a_n56_158# Gnd nfet w=4 l=3
+ ad=0 pd=0 as=0 ps=0 
C0 myVdd myClr 2.7fF
C1 myVdd myD 2.7fF
C2 myVdd not_0/myOut 2.2fF
C3 myGnd dff1_0/not_0/myA 5.9fF
C4 myGnd dff1_0/a_n56_158# 2.2fF
C5 myVdd myOut2 3.6fF
C6 myVdd dff1_0/not_0/myA 5.6fF
C7 myVdd dff1_0/not_2/myA 2.5fF
C8 myVdd myGnd 11.4fF
C9 myGnd dff1_0/gate_1/myD 2.9fF
C10 myOut2 gnd! 58.2fF
C11 dff1_0/a_n56_158# gnd! 23.9fF
C12 dff1_0/a_n81_156# gnd! 25.2fF
C13 myOut1 gnd! 74.5fF
C14 dff1_0/a_n133_170# gnd! 25.2fF
C15 myClr gnd! 14.9fF
C16 dff1_0/clr_0/a_33_50# gnd! 25.2fF
C17 myD gnd! 36.5fF
C18 dff1_0/clr_0/a_n13_27# gnd! 23.5fF
C19 dff1_0/gate_0/myC gnd! 42.5fF
C20 dff1_0/gate_0/myD gnd! 17.8fF
C21 dff1_0/gate_0/a_3_46# gnd! 25.2fF
C22 dff1_0/not_0/myA gnd! 246.4fF
C23 dff1_0/gate_1/a_3_46# gnd! 25.2fF
C24 dff1_0/not_1/myA gnd! 43.3fF
C25 dff1_0/gate_1/myD gnd! 23.9fF
C26 dff1_0/not_2/myA gnd! 48.7fF
C27 dff1_0/not_4/myOut gnd! 32.8fF
C28 not_0/myOut gnd! 25.7fF
C29 myGnd gnd! 249.2fF
C30 not_0/myA gnd! 16.0fF
C31 myVdd gnd! 467.0fF
C32 myClk gnd! 13.3fF

.include ../usc-spice.usc-spice

Vgnd1 myGnd 0 DC 0V
Vgnd2 gnd! 0 DC 0V

VVdd myVdd 0 DC 2.8V

Vin1 myD 0 pulse(0 2.8v 0ns 0.1ns 0.1ns 100ns 200ns)
Vin2 myClk 0 pulse(0 2.8v 0ns 0.1ns 0.1ns 32ns 64ns)
Vin3 myClr 0 pulse(0 2.8v 0ns 0.1ns 0.1ns 250ns 500ns)

.tran 1ns 1400ns
.probe
.control
run
plot myClk myD+4 myClr+8 myOut2+12 myOut1+16
.endc
.end