* SPICE3 file created from xor.ext - technology: scmos

.option scale=1u

M1000 a_n9_n15# myIna myVdd w_n26_n2# pfet w=6 l=4
+ ad=42 pd=26 as=189 ps=96 
M1001 a_23_n15# myInb myVdd w_n26_n2# pfet w=6 l=4
+ ad=42 pd=26 as=0 ps=0 
M1002 a_n9_n15# myIna myGnd Gnd nfet w=6 l=4
+ ad=48 pd=28 as=252 ps=132 
M1003 a_23_n15# myInb myGnd Gnd nfet w=6 l=4
+ ad=48 pd=28 as=0 ps=0 
M1004 a_n9_n38# myIna myGnd Gnd nfet w=6 l=4
+ ad=162 pd=78 as=0 ps=0 
M1005 myOut a_n9_n15# a_n9_n38# Gnd nfet w=6 l=4
+ ad=72 pd=36 as=0 ps=0 
M1006 a_n9_n38# myInb myOut Gnd nfet w=6 l=4
+ ad=0 pd=0 as=0 ps=0 
M1007 myGnd a_23_n15# a_n9_n38# Gnd nfet w=6 l=4
+ ad=0 pd=0 as=0 ps=0 
M1008 myOut myIna a_n32_n57# w_n33_n60# pfet w=7 l=4
+ ad=84 pd=38 as=217 ps=90 
M1009 a_7_n57# a_n9_n15# myOut w_n33_n60# pfet w=7 l=4
+ ad=84 pd=38 as=0 ps=0 
M1010 myVdd myInb a_7_n57# w_n33_n60# pfet w=7 l=4
+ ad=0 pd=0 as=0 ps=0 
M1011 a_n32_n57# a_23_n15# myVdd w_n33_n60# pfet w=7 l=4
+ ad=0 pd=0 as=0 ps=0 
C0 a_n32_n57# gnd! 12.0fF
C1 myOut gnd! 8.1fF
C2 a_n9_n38# gnd! 5.0fF
C3 myGnd gnd! 21.4fF
C4 a_23_n15# gnd! 18.2fF
C5 a_n9_n15# gnd! 17.2fF
C6 myVdd gnd! 40.3fF
C7 myInb gnd! 18.4fF
C8 myIna gnd! 18.4fF

.include ../usc-spice.usc-spice

Vgnd1 myGnd 0 DC 0V
Vgnd2 gnd! 0 DC 0V

VVdd myVdd 0 DC 2.8V

Vin1 myIna 0 pulse(0 2.8v 0ns 0.1ns 0.1ns 64ns 128ns)
Vin2 myInb 0 pulse(0 2.8v 0ns 0.1ns 0.1ns 128ns 256ns)

.tran 1ns 1000ns
.probe
.control
run
plot myIna myInb+4 myOut+8
.endc
.end

