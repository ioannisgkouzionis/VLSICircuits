magic
tech scmos
timestamp 1477328863
<< nwell >>
rect -48 110 42 120
rect 69 110 159 120
rect -27 44 35 54
rect 76 44 138 54
<< polysilicon >>
rect -33 117 -29 125
rect -14 117 -10 125
rect 2 117 6 125
rect 18 117 22 125
rect 89 117 93 125
rect 105 117 109 125
rect 121 117 125 125
rect 140 117 144 125
rect -33 90 -29 110
rect -14 90 -10 110
rect 2 90 6 110
rect 18 90 22 110
rect 89 98 93 110
rect 89 90 93 93
rect 105 90 109 110
rect 121 90 125 110
rect 140 90 144 110
rect -33 65 -29 84
rect -14 67 -10 84
rect 2 65 6 84
rect 18 67 22 84
rect 89 67 93 84
rect 105 65 109 84
rect 121 67 125 84
rect 140 65 144 84
rect -14 51 -10 61
rect 18 51 22 61
rect 89 51 93 61
rect 121 51 125 61
rect -14 34 -10 45
rect 18 35 22 45
rect 89 43 93 45
rect 121 31 125 45
rect 9 -1 25 1
rect 30 -1 67 1
rect 9 -2 67 -1
rect 9 -11 12 -2
rect 24 -11 27 -9
rect 42 -11 46 -9
rect 64 -11 67 -2
rect 73 -11 77 -1
rect 115 -11 119 -7
rect 9 -35 12 -18
rect 24 -35 27 -18
rect 42 -35 46 -18
rect 64 -35 67 -18
rect 73 -35 77 -18
rect 115 -24 119 -18
rect 117 -30 119 -24
rect 115 -34 119 -30
rect 9 -45 12 -42
rect 24 -47 27 -42
rect 42 -45 46 -42
rect 64 -45 67 -42
rect 73 -47 77 -42
rect 115 -45 119 -41
rect 24 -49 77 -47
<< ndiffusion >>
rect -45 89 -33 90
rect -45 85 -44 89
rect -40 85 -33 89
rect -45 84 -33 85
rect -29 89 -14 90
rect -29 85 -24 89
rect -20 85 -14 89
rect -29 84 -14 85
rect -10 89 2 90
rect -10 85 -6 89
rect -2 85 2 89
rect -10 84 2 85
rect 6 89 18 90
rect 6 85 10 89
rect 14 85 18 89
rect 6 84 18 85
rect 22 89 39 90
rect 22 85 24 89
rect 28 85 39 89
rect 22 84 39 85
rect 72 89 89 90
rect 72 85 83 89
rect 87 85 89 89
rect 72 84 89 85
rect 93 89 105 90
rect 93 85 97 89
rect 101 85 105 89
rect 93 84 105 85
rect 109 89 121 90
rect 109 85 113 89
rect 117 85 121 89
rect 109 84 121 85
rect 125 89 140 90
rect 125 85 131 89
rect 135 85 140 89
rect 125 84 140 85
rect 144 89 156 90
rect 144 85 151 89
rect 155 85 156 89
rect 144 84 156 85
rect -22 66 -14 67
rect -22 62 -20 66
rect -16 62 -14 66
rect -22 61 -14 62
rect -10 66 -4 67
rect -10 62 -9 66
rect -5 62 -4 66
rect -10 61 -4 62
rect 10 66 18 67
rect 10 62 12 66
rect 16 62 18 66
rect 10 61 18 62
rect 22 66 29 67
rect 22 62 24 66
rect 28 62 29 66
rect 22 61 29 62
rect 82 66 89 67
rect 82 62 83 66
rect 87 62 89 66
rect 82 61 89 62
rect 93 66 101 67
rect 93 62 95 66
rect 99 62 101 66
rect 93 61 101 62
rect 115 66 121 67
rect 115 62 116 66
rect 120 62 121 66
rect 115 61 121 62
rect 125 66 133 67
rect 125 62 127 66
rect 131 62 133 66
rect 125 61 133 62
rect 105 -35 115 -34
rect -1 -36 9 -35
rect -1 -41 1 -36
rect 6 -41 9 -36
rect -1 -42 9 -41
rect 12 -36 24 -35
rect 12 -41 16 -36
rect 21 -41 24 -36
rect 12 -42 24 -41
rect 27 -36 42 -35
rect 27 -41 31 -36
rect 36 -41 42 -36
rect 27 -42 42 -41
rect 46 -36 64 -35
rect 46 -41 53 -36
rect 58 -41 64 -36
rect 46 -42 64 -41
rect 67 -42 73 -35
rect 77 -36 90 -35
rect 77 -41 81 -36
rect 86 -41 90 -36
rect 105 -40 107 -35
rect 112 -40 115 -35
rect 105 -41 115 -40
rect 119 -35 130 -34
rect 119 -40 123 -35
rect 128 -40 130 -35
rect 119 -41 130 -40
rect 77 -42 90 -41
<< pdiffusion >>
rect -45 116 -33 117
rect -45 112 -44 116
rect -40 112 -33 116
rect -45 110 -33 112
rect -29 116 -14 117
rect -29 112 -24 116
rect -20 112 -14 116
rect -29 110 -14 112
rect -10 110 2 117
rect 6 116 18 117
rect 6 112 9 116
rect 13 112 18 116
rect 6 110 18 112
rect 22 116 41 117
rect 22 112 24 116
rect 28 112 41 116
rect 22 110 41 112
rect 70 116 89 117
rect 70 112 83 116
rect 87 112 89 116
rect 70 110 89 112
rect 93 116 105 117
rect 93 112 98 116
rect 102 112 105 116
rect 93 110 105 112
rect 109 110 121 117
rect 125 116 140 117
rect 125 112 131 116
rect 135 112 140 116
rect 125 110 140 112
rect 144 116 156 117
rect 144 112 151 116
rect 155 112 156 116
rect 144 110 156 112
rect -21 50 -14 51
rect -21 46 -20 50
rect -16 46 -14 50
rect -21 45 -14 46
rect -10 50 -3 51
rect -10 46 -8 50
rect -4 46 -3 50
rect -10 45 -3 46
rect 11 50 18 51
rect 11 46 12 50
rect 16 46 18 50
rect 11 45 18 46
rect 22 50 29 51
rect 22 46 24 50
rect 28 46 29 50
rect 22 45 29 46
rect 82 50 89 51
rect 82 46 83 50
rect 87 46 89 50
rect 82 45 89 46
rect 93 50 100 51
rect 93 46 95 50
rect 99 46 100 50
rect 93 45 100 46
rect 114 50 121 51
rect 114 46 115 50
rect 119 46 121 50
rect 114 45 121 46
rect 125 50 132 51
rect 125 46 127 50
rect 131 46 132 50
rect 125 45 132 46
rect -1 -12 9 -11
rect -1 -17 1 -12
rect 6 -17 9 -12
rect -1 -18 9 -17
rect 12 -12 24 -11
rect 12 -17 15 -12
rect 20 -17 24 -12
rect 12 -18 24 -17
rect 27 -12 42 -11
rect 27 -17 31 -12
rect 36 -17 42 -12
rect 27 -18 42 -17
rect 46 -12 64 -11
rect 46 -17 52 -12
rect 57 -17 64 -12
rect 46 -18 64 -17
rect 67 -18 73 -11
rect 77 -12 89 -11
rect 77 -17 81 -12
rect 86 -17 89 -12
rect 77 -18 89 -17
rect 105 -12 115 -11
rect 105 -17 107 -12
rect 112 -17 115 -12
rect 105 -18 115 -17
rect 119 -12 130 -11
rect 119 -17 123 -12
rect 128 -17 130 -12
rect 119 -18 130 -17
<< metal1 >>
rect 62 140 220 145
rect -44 125 28 128
rect -44 116 -40 125
rect 24 116 28 125
rect -24 109 -20 112
rect -61 106 -20 109
rect -61 43 -57 106
rect 9 98 13 112
rect 62 109 66 140
rect 83 125 155 128
rect 83 116 87 125
rect 151 116 155 125
rect 98 109 102 112
rect 131 109 135 112
rect 62 106 117 109
rect 131 106 172 109
rect -6 93 89 98
rect -6 89 -2 93
rect 113 89 117 106
rect -44 74 -40 85
rect -24 82 -20 85
rect 10 82 14 85
rect -24 79 14 82
rect 24 74 28 85
rect 83 74 87 85
rect 97 82 101 85
rect 131 82 135 85
rect 97 79 135 82
rect 151 74 155 85
rect -44 69 153 74
rect -9 66 -5 69
rect 24 66 28 69
rect -33 58 -29 61
rect -20 58 -16 62
rect -33 54 -16 58
rect 2 58 6 61
rect 83 66 87 69
rect 116 66 120 69
rect 12 58 16 62
rect 2 55 16 58
rect -20 50 -16 54
rect 12 50 16 55
rect 95 58 99 62
rect 105 58 109 61
rect 95 55 109 58
rect 127 58 131 62
rect 140 58 144 61
rect 95 50 99 55
rect 127 54 144 58
rect 127 50 131 54
rect -8 43 -4 46
rect 24 43 28 46
rect 83 43 87 46
rect 115 43 119 46
rect 168 43 172 106
rect -61 38 172 43
rect -61 20 -57 38
rect -30 28 -14 34
rect -14 27 -10 28
rect 22 31 40 35
rect 18 30 22 31
rect 64 26 121 31
rect -73 17 57 20
rect 25 3 30 5
rect 42 -5 46 2
rect 1 -9 36 -6
rect 52 -6 57 17
rect 73 3 77 26
rect 52 -9 112 -6
rect 1 -12 6 -9
rect 31 -12 36 -9
rect 52 -12 57 -9
rect 107 -12 112 -9
rect 15 -20 20 -17
rect 81 -20 86 -17
rect 15 -23 86 -20
rect 81 -24 86 -23
rect 123 -23 128 -17
rect 81 -30 113 -24
rect 123 -28 217 -23
rect 16 -33 86 -30
rect 16 -36 21 -33
rect 81 -36 86 -33
rect 123 -35 128 -28
rect 1 -51 6 -41
rect 31 -51 36 -41
rect 1 -54 36 -51
rect 53 -51 58 -41
rect 107 -51 112 -40
rect 53 -56 112 -51
rect 53 -60 58 -56
rect -70 -67 94 -60
<< metal2 >>
rect 159 69 199 74
rect -14 27 -10 28
rect -14 9 -10 23
rect 18 18 22 26
rect 18 15 46 18
rect -14 5 25 9
rect 42 6 46 15
rect 191 -60 199 69
rect 103 -67 199 -60
<< ntransistor >>
rect -33 84 -29 90
rect -14 84 -10 90
rect 2 84 6 90
rect 18 84 22 90
rect 89 84 93 90
rect 105 84 109 90
rect 121 84 125 90
rect 140 84 144 90
rect -14 61 -10 67
rect 18 61 22 67
rect 89 61 93 67
rect 121 61 125 67
rect 9 -42 12 -35
rect 24 -42 27 -35
rect 42 -42 46 -35
rect 64 -42 67 -35
rect 73 -42 77 -35
rect 115 -41 119 -34
<< ptransistor >>
rect -33 110 -29 117
rect -14 110 -10 117
rect 2 110 6 117
rect 18 110 22 117
rect 89 110 93 117
rect 105 110 109 117
rect 121 110 125 117
rect 140 110 144 117
rect -14 45 -10 51
rect 18 45 22 51
rect 89 45 93 51
rect 121 45 125 51
rect 9 -18 12 -11
rect 24 -18 27 -11
rect 42 -18 46 -11
rect 64 -18 67 -11
rect 73 -18 77 -11
rect 115 -18 119 -11
<< polycontact >>
rect 89 93 93 98
rect -33 61 -29 65
rect 2 61 6 65
rect 105 61 109 65
rect 140 61 144 65
rect -14 28 -10 34
rect 18 31 22 35
rect 121 26 125 31
rect 25 -1 30 3
rect 42 -9 46 -5
rect 73 -1 77 3
rect 113 -30 117 -24
<< ndcontact >>
rect -44 85 -40 89
rect -24 85 -20 89
rect -6 85 -2 89
rect 10 85 14 89
rect 24 85 28 89
rect 83 85 87 89
rect 97 85 101 89
rect 113 85 117 89
rect 131 85 135 89
rect 151 85 155 89
rect -20 62 -16 66
rect -9 62 -5 66
rect 12 62 16 66
rect 24 62 28 66
rect 83 62 87 66
rect 95 62 99 66
rect 116 62 120 66
rect 127 62 131 66
rect 1 -41 6 -36
rect 16 -41 21 -36
rect 31 -41 36 -36
rect 53 -41 58 -36
rect 81 -41 86 -36
rect 107 -40 112 -35
rect 123 -40 128 -35
<< pdcontact >>
rect -44 112 -40 116
rect -24 112 -20 116
rect 9 112 13 116
rect 24 112 28 116
rect 83 112 87 116
rect 98 112 102 116
rect 131 112 135 116
rect 151 112 155 116
rect -20 46 -16 50
rect -8 46 -4 50
rect 12 46 16 50
rect 24 46 28 50
rect 83 46 87 50
rect 95 46 99 50
rect 115 46 119 50
rect 127 46 131 50
rect 1 -17 6 -12
rect 15 -17 20 -12
rect 31 -17 36 -12
rect 52 -17 57 -12
rect 81 -17 86 -12
rect 107 -17 112 -12
rect 123 -17 128 -12
<< m2contact >>
rect 153 69 159 74
rect -14 23 -10 27
rect 18 26 22 30
rect 25 5 30 9
rect 42 2 46 6
rect 94 -67 103 -60
<< labels >>
rlabel metal1 -71 18 -71 18 3 myVdd
rlabel metal1 38 33 38 33 1 myA
rlabel metal1 -26 30 -26 30 1 myB
rlabel metal1 -65 -63 -65 -63 1 myGnd
rlabel metal1 68 28 68 28 1 myCin
rlabel metal1 211 -26 211 -26 1 myCout
rlabel metal1 216 143 216 143 6 mySum
<< end >>
