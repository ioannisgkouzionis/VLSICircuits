magic
tech scmos
timestamp 1478865149
<< polysilicon >>
rect -133 181 -108 184
rect -133 177 -130 181
rect -133 170 -130 172
rect -133 162 -130 166
rect -112 161 -108 181
rect -133 148 -130 158
rect -81 181 -56 184
rect -81 161 -77 181
rect -59 177 -56 181
rect 3 178 6 182
rect -59 170 -56 172
rect 3 169 6 173
rect -59 162 -56 166
rect 5 165 6 169
rect 3 160 6 165
rect -59 148 -56 158
rect 3 152 6 156
rect -133 139 -130 143
rect -131 135 -130 139
rect -133 130 -130 135
rect -59 139 -56 143
rect -59 135 -58 139
rect 4 136 7 140
rect -59 130 -56 135
rect 4 127 7 131
rect -133 122 -130 126
rect -59 122 -56 126
rect 4 123 5 127
rect 4 118 7 123
rect 4 110 7 114
<< ndiffusion >>
rect -145 158 -142 162
rect -138 158 -133 162
rect -130 158 -123 162
rect -119 158 -117 162
rect -72 158 -70 162
rect -66 158 -59 162
rect -56 158 -51 162
rect -47 158 -44 162
rect -8 156 -5 160
rect -1 156 3 160
rect 6 156 12 160
rect 16 156 18 160
rect -144 126 -141 130
rect -137 126 -133 130
rect -130 126 -124 130
rect -120 126 -118 130
rect -71 126 -69 130
rect -65 126 -59 130
rect -56 126 -52 130
rect -48 126 -45 130
rect -8 114 -6 118
rect -2 114 4 118
rect 7 114 11 118
rect 15 114 18 118
<< pdiffusion >>
rect -144 173 -142 177
rect -138 173 -133 177
rect -144 172 -133 173
rect -130 173 -123 177
rect -119 173 -118 177
rect -130 172 -118 173
rect -71 173 -70 177
rect -66 173 -59 177
rect -71 172 -59 173
rect -56 173 -51 177
rect -47 173 -45 177
rect -9 174 -7 178
rect -3 174 3 178
rect -9 173 3 174
rect 6 174 12 178
rect 16 174 17 178
rect 6 173 17 174
rect -56 172 -45 173
rect -145 144 -143 148
rect -139 144 -133 148
rect -145 143 -133 144
rect -130 144 -124 148
rect -120 144 -119 148
rect -130 143 -119 144
rect -70 144 -69 148
rect -65 144 -59 148
rect -70 143 -59 144
rect -56 144 -50 148
rect -46 144 -44 148
rect -56 143 -44 144
rect -7 132 -6 136
rect -2 132 4 136
rect -7 131 4 132
rect 7 132 13 136
rect 17 132 19 136
rect 7 131 19 132
<< metal1 >>
rect -80 208 -70 214
rect -530 198 -352 200
rect -268 202 -220 206
rect -530 194 -346 198
rect -530 36 -520 194
rect -448 188 -440 194
rect -350 188 -346 194
rect -312 194 -234 198
rect -312 170 -308 194
rect -240 170 -234 194
rect -224 184 -218 202
rect -78 198 -74 208
rect -96 194 -18 198
rect -194 170 -180 172
rect -388 164 -366 170
rect -318 166 -304 170
rect -256 164 -246 170
rect -240 164 -224 170
rect -194 169 -150 170
rect -142 169 -138 173
rect -194 165 -138 169
rect -194 164 -146 165
rect -513 156 -500 160
rect -376 134 -362 140
rect -470 104 -464 117
rect -376 62 -370 134
rect -358 104 -352 122
rect -358 92 -352 98
rect -268 94 -264 124
rect -358 88 -268 92
rect -346 78 -340 88
rect -376 58 -368 62
rect -336 58 -314 64
rect -320 54 -314 58
rect -260 54 -256 140
rect -250 130 -246 164
rect -238 148 -216 150
rect -232 144 -216 148
rect -250 122 -230 130
rect -188 128 -180 164
rect -142 162 -138 165
rect -133 154 -130 186
rect -123 170 -119 173
rect -96 170 -92 194
rect -70 170 -66 173
rect -123 166 -66 170
rect -123 162 -119 166
rect -70 162 -66 166
rect -143 151 -130 154
rect -143 148 -139 151
rect -148 140 -141 141
rect -194 122 -180 128
rect -160 139 -141 140
rect -124 140 -120 144
rect -112 140 -108 156
rect -160 135 -135 139
rect -124 136 -108 140
rect -81 140 -77 156
rect -59 154 -56 186
rect -51 169 -47 173
rect -24 170 -18 194
rect -7 178 -3 184
rect 12 170 16 174
rect 22 170 64 172
rect -40 169 -30 170
rect -51 165 -30 169
rect -51 162 -47 165
rect -40 164 -30 165
rect -24 169 -8 170
rect -24 165 1 169
rect 12 165 64 170
rect -24 164 -8 165
rect 12 164 58 165
rect -59 151 -46 154
rect -50 148 -46 151
rect -69 140 -65 144
rect -81 136 -65 140
rect -44 139 -40 140
rect -160 134 -146 135
rect -206 94 -200 108
rect -160 54 -154 134
rect -124 130 -120 136
rect -69 130 -65 136
rect -54 135 -40 139
rect -141 125 -137 126
rect -141 120 -136 125
rect -142 94 -136 120
rect -52 108 -48 126
rect -52 94 -48 104
rect -44 104 -40 135
rect -34 130 -30 164
rect 12 160 16 164
rect -5 152 -1 156
rect 13 136 17 140
rect -34 128 -14 130
rect -6 128 -2 132
rect 28 128 36 164
rect -34 124 -2 128
rect 22 127 36 128
rect -34 122 -14 124
rect -6 118 -2 124
rect 9 123 36 127
rect 22 122 36 123
rect 11 112 15 114
rect -44 100 6 104
rect -136 92 -48 94
rect -136 88 -54 92
rect -66 68 -10 78
rect 2 54 8 68
rect 22 64 26 76
rect -320 46 58 54
rect 92 46 110 52
rect -346 36 -336 44
rect -530 26 -336 36
<< metal2 >>
rect -346 202 -274 206
rect -214 202 -174 206
rect -346 200 -270 202
rect -276 190 -270 200
rect -178 190 -174 202
rect -178 186 -134 190
rect -130 186 -60 190
rect -56 186 -8 190
rect -178 150 -174 186
rect -2 186 44 190
rect -240 144 -238 148
rect -512 128 -502 134
rect -464 98 -358 104
rect -240 94 -232 144
rect -204 146 -174 150
rect -22 148 -6 152
rect -204 144 -198 146
rect -22 108 -16 148
rect 38 146 44 186
rect 38 144 88 146
rect 18 140 88 144
rect -48 106 10 108
rect -48 104 16 106
rect -264 88 -206 94
rect -200 88 -142 94
rect -78 6 -68 68
rect -54 64 -48 88
rect 82 82 88 140
rect 82 78 136 82
rect 82 70 88 78
rect -54 60 22 64
rect 20 28 26 60
rect 80 28 86 32
rect 20 20 86 28
rect 124 6 136 78
rect -78 -4 136 6
<< ntransistor >>
rect -133 158 -130 162
rect -59 158 -56 162
rect 3 156 6 160
rect -133 126 -130 130
rect -59 126 -56 130
rect 4 114 7 118
<< ptransistor >>
rect -133 172 -130 177
rect -59 172 -56 177
rect 3 173 6 178
rect -133 143 -130 148
rect -59 143 -56 148
rect 4 131 7 136
<< polycontact >>
rect -112 156 -108 161
rect 1 165 5 169
rect -81 156 -77 161
rect -135 135 -131 139
rect -58 135 -54 139
rect 5 123 9 127
<< ndcontact >>
rect -142 158 -138 162
rect -123 158 -119 162
rect -70 158 -66 162
rect -51 158 -47 162
rect -5 156 -1 160
rect 12 156 16 160
rect -141 126 -137 130
rect -124 126 -120 130
rect -69 126 -65 130
rect -52 126 -48 130
rect -6 114 -2 118
rect 11 114 15 118
<< pdcontact >>
rect -142 173 -138 177
rect -123 173 -119 177
rect -70 173 -66 177
rect -51 173 -47 177
rect -7 174 -3 178
rect 12 174 16 178
rect -143 144 -139 148
rect -124 144 -120 148
rect -69 144 -65 148
rect -50 144 -46 148
rect -6 132 -2 136
rect 13 132 17 136
<< m2contact >>
rect -352 198 -346 206
rect -274 202 -268 206
rect -220 202 -214 206
rect -276 186 -270 190
rect -134 186 -130 190
rect -470 98 -464 104
rect -358 98 -352 104
rect -268 88 -264 94
rect -238 144 -232 148
rect -204 140 -198 144
rect -60 186 -56 190
rect -8 184 -2 190
rect -206 88 -200 94
rect -52 104 -48 108
rect -6 148 0 152
rect 12 140 18 144
rect 10 106 16 112
rect -142 88 -136 94
rect -54 88 -48 92
rect -78 68 -66 78
rect 82 64 88 70
rect 22 60 26 64
rect 80 32 86 36
use clr  clr_0
timestamp 1478860239
transform 1 0 -470 0 1 120
box -36 -4 83 70
use gate  gate_0
timestamp 1478855084
transform 1 0 -352 0 1 124
box -16 -4 35 64
use gate  gate_1
timestamp 1478855084
transform -1 0 -269 0 1 124
box -16 -4 35 64
use not  not_1
timestamp 1478778185
transform 1 0 -199 0 1 167
box -29 -17 7 17
use not  not_2
timestamp 1478778185
transform -1 0 -223 0 1 125
box -29 -17 7 17
use not  not_0
timestamp 1478778185
transform -1 0 -363 0 -1 61
box -29 -17 7 17
use not  not_4
timestamp 1478778185
transform 0 -1 5 1 0 95
box -29 -17 7 17
use not  not_3
timestamp 1478778185
transform -1 0 63 0 1 49
box -29 -17 7 17
<< labels >>
rlabel metal1 -510 158 -510 158 3 myClr
rlabel metal2 -508 132 -508 132 3 myD
rlabel metal1 108 48 108 48 7 myClk
rlabel metal1 -382 197 -382 197 1 myVdd
rlabel metal2 -437 99 -437 99 1 myGnd
rlabel metal1 -75 211 -75 211 5 myOut1
rlabel metal1 60 166 60 166 1 myOut2
<< end >>
