magic
tech scmos
timestamp 1478778185
<< polysilicon >>
rect -14 11 -11 15
rect -14 2 -11 6
rect -12 -2 -11 2
rect -14 -7 -11 -2
rect -14 -15 -11 -11
<< ndiffusion >>
rect -25 -11 -22 -7
rect -18 -11 -14 -7
rect -11 -11 -5 -7
rect -1 -11 1 -7
<< pdiffusion >>
rect -26 7 -24 11
rect -20 7 -14 11
rect -26 6 -14 7
rect -11 7 -5 11
rect -1 7 0 11
rect -11 6 0 7
<< metal1 >>
rect -24 11 -20 17
rect -5 3 -1 7
rect -29 -2 -16 2
rect -5 -1 7 3
rect -5 -7 -1 -1
rect -22 -17 -18 -11
<< ntransistor >>
rect -14 -11 -11 -7
<< ptransistor >>
rect -14 6 -11 11
<< polycontact >>
rect -16 -2 -12 2
<< ndcontact >>
rect -22 -11 -18 -7
rect -5 -11 -1 -7
<< pdcontact >>
rect -24 7 -20 11
rect -5 7 -1 11
<< labels >>
rlabel metal1 -22 15 -22 15 5 myVdd
rlabel metal1 -27 0 -27 0 3 myA
rlabel metal1 5 0 5 0 7 myOut
rlabel metal1 -20 -15 -20 -15 1 myGnd
<< end >>
