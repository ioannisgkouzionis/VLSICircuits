magic
tech scmos
timestamp 1479555546
<< polysilicon >>
rect 27 156 29 167
rect 57 156 59 167
rect 27 139 29 150
rect 57 139 59 150
rect 15 121 17 136
rect 27 121 29 136
rect 45 121 47 136
rect 15 107 17 118
rect 27 107 29 118
rect 57 121 59 136
rect 104 130 138 132
rect 94 126 96 128
rect 104 126 106 130
rect 116 126 118 128
rect 129 126 131 128
rect 136 126 138 130
rect 154 126 156 128
rect 45 107 47 118
rect 57 107 59 118
rect 94 113 96 123
rect 104 113 106 123
rect 116 113 118 123
rect 129 113 131 123
rect 136 113 138 123
rect 154 113 156 123
rect 15 99 17 101
rect 27 99 29 101
rect 45 99 47 101
rect 57 99 59 101
rect 94 99 96 107
rect 104 105 106 107
rect 116 106 118 107
rect 129 99 131 107
rect 136 99 138 107
rect 154 105 156 107
rect 86 95 92 97
rect 96 97 131 99
rect 86 75 88 95
rect 111 91 128 93
rect 116 75 118 83
rect 143 75 145 77
rect 173 75 175 83
rect 86 58 88 69
rect 116 58 118 69
rect 143 58 145 69
rect 173 58 175 69
rect 74 40 76 55
rect 86 40 88 55
rect 104 40 106 55
rect 74 26 76 37
rect 86 26 88 37
rect 116 40 118 55
rect 143 40 145 55
rect 155 40 157 55
rect 173 40 175 55
rect 104 26 106 37
rect 116 26 118 37
rect 143 34 145 37
rect 143 22 145 30
rect 155 22 157 37
rect 185 40 187 55
rect 173 22 175 37
rect 185 22 187 37
rect 74 18 76 20
rect 86 18 88 20
rect 104 18 106 20
rect 116 18 118 20
rect 143 14 145 16
rect 155 14 157 16
rect 173 14 175 16
rect 185 14 187 16
<< ndiffusion >>
rect 18 136 20 139
rect 24 136 27 139
rect 29 136 32 139
rect 36 136 38 139
rect 48 136 50 139
rect 54 136 57 139
rect 59 136 62 139
rect 66 136 68 139
rect 6 118 8 121
rect 12 118 15 121
rect 17 118 20 121
rect 24 118 27 121
rect 29 118 35 121
rect 39 118 45 121
rect 47 118 50 121
rect 87 123 88 126
rect 92 123 94 126
rect 96 123 98 126
rect 102 123 104 126
rect 106 123 108 126
rect 112 123 116 126
rect 118 123 122 126
rect 126 123 129 126
rect 131 123 136 126
rect 138 123 140 126
rect 144 123 145 126
rect 148 123 149 126
rect 153 123 154 126
rect 156 123 157 126
rect 161 123 163 126
rect 54 118 57 121
rect 59 118 62 121
rect 66 118 68 121
rect 77 55 79 58
rect 83 55 86 58
rect 88 55 91 58
rect 95 55 97 58
rect 107 55 109 58
rect 113 55 116 58
rect 118 55 121 58
rect 125 55 127 58
rect 134 55 136 58
rect 140 55 143 58
rect 145 55 148 58
rect 152 55 154 58
rect 164 55 166 58
rect 170 55 173 58
rect 175 55 178 58
rect 182 55 184 58
rect 65 37 67 40
rect 71 37 74 40
rect 76 37 79 40
rect 83 37 86 40
rect 88 37 94 40
rect 98 37 104 40
rect 106 37 109 40
rect 113 37 116 40
rect 118 37 121 40
rect 125 37 127 40
rect 134 37 136 40
rect 140 37 143 40
rect 145 37 148 40
rect 152 37 155 40
rect 157 37 163 40
rect 167 37 173 40
rect 175 37 178 40
rect 182 37 185 40
rect 187 37 190 40
rect 194 37 196 40
<< pdiffusion >>
rect 18 155 27 156
rect 18 151 20 155
rect 24 151 27 155
rect 18 150 27 151
rect 29 155 38 156
rect 29 151 32 155
rect 36 151 38 155
rect 29 150 38 151
rect 48 155 57 156
rect 48 151 50 155
rect 54 151 57 155
rect 48 150 57 151
rect 59 155 68 156
rect 59 151 62 155
rect 66 151 68 155
rect 59 150 68 151
rect 87 112 94 113
rect 87 108 88 112
rect 92 108 94 112
rect 87 107 94 108
rect 96 112 104 113
rect 96 108 98 112
rect 102 108 104 112
rect 96 107 104 108
rect 106 112 116 113
rect 106 108 108 112
rect 112 108 116 112
rect 106 107 116 108
rect 118 112 129 113
rect 118 108 122 112
rect 126 108 129 112
rect 118 107 129 108
rect 131 107 136 113
rect 138 112 145 113
rect 138 108 140 112
rect 144 108 145 112
rect 138 107 145 108
rect 148 112 154 113
rect 148 108 149 112
rect 153 108 154 112
rect 148 107 154 108
rect 156 112 163 113
rect 156 108 157 112
rect 161 108 163 112
rect 156 107 163 108
rect 6 106 15 107
rect 6 102 8 106
rect 12 102 15 106
rect 6 101 15 102
rect 17 106 27 107
rect 17 102 20 106
rect 24 102 27 106
rect 17 101 27 102
rect 29 101 45 107
rect 47 106 57 107
rect 47 102 50 106
rect 54 102 57 106
rect 47 101 57 102
rect 59 106 68 107
rect 59 102 62 106
rect 66 102 68 106
rect 59 101 68 102
rect 77 74 86 75
rect 77 70 79 74
rect 83 70 86 74
rect 77 69 86 70
rect 88 74 97 75
rect 88 70 91 74
rect 95 70 97 74
rect 88 69 97 70
rect 107 74 116 75
rect 107 70 109 74
rect 113 70 116 74
rect 107 69 116 70
rect 118 74 127 75
rect 118 70 121 74
rect 125 70 127 74
rect 118 69 127 70
rect 134 74 143 75
rect 134 70 136 74
rect 140 70 143 74
rect 134 69 143 70
rect 145 74 154 75
rect 145 70 148 74
rect 152 70 154 74
rect 145 69 154 70
rect 164 74 173 75
rect 164 70 166 74
rect 170 70 173 74
rect 164 69 173 70
rect 175 74 184 75
rect 175 70 178 74
rect 182 70 184 74
rect 175 69 184 70
rect 65 25 74 26
rect 65 21 67 25
rect 71 21 74 25
rect 65 20 74 21
rect 76 25 86 26
rect 76 21 79 25
rect 83 21 86 25
rect 76 20 86 21
rect 88 20 104 26
rect 106 25 116 26
rect 106 21 109 25
rect 113 21 116 25
rect 106 20 116 21
rect 118 25 127 26
rect 118 21 121 25
rect 125 21 127 25
rect 118 20 127 21
rect 134 21 143 22
rect 134 17 136 21
rect 140 17 143 21
rect 134 16 143 17
rect 145 21 155 22
rect 145 17 148 21
rect 152 17 155 21
rect 145 16 155 17
rect 157 16 173 22
rect 175 21 185 22
rect 175 17 178 21
rect 182 17 185 21
rect 175 16 185 17
rect 187 21 196 22
rect 187 17 190 21
rect 194 17 196 21
rect 187 16 196 17
<< metal1 >>
rect 2 158 74 161
rect 2 112 5 158
rect 32 155 35 158
rect 62 155 65 158
rect 20 146 23 151
rect 50 146 53 151
rect 14 143 23 146
rect 14 140 17 143
rect 20 140 23 143
rect 44 143 53 146
rect 44 140 47 143
rect 50 140 53 143
rect 71 141 74 158
rect 71 137 121 141
rect 32 133 35 136
rect 62 133 65 136
rect 9 130 70 133
rect 9 122 12 130
rect 21 124 53 127
rect 21 122 24 124
rect 50 122 53 124
rect 62 122 65 130
rect 89 130 111 133
rect 89 127 92 130
rect 108 127 111 130
rect 122 130 144 133
rect 148 130 152 133
rect 122 127 125 130
rect 149 127 152 130
rect 99 119 102 123
rect 140 119 143 123
rect 158 119 161 123
rect 36 112 39 117
rect 99 116 150 119
rect 99 112 102 116
rect 140 112 143 116
rect 158 116 167 119
rect 158 112 161 116
rect 2 109 23 112
rect 36 109 82 112
rect 20 106 23 109
rect 51 106 54 109
rect 9 99 12 102
rect 62 99 65 102
rect 9 96 65 99
rect 79 99 82 109
rect 89 105 92 108
rect 108 105 111 108
rect 89 102 111 105
rect 122 105 125 108
rect 149 105 152 108
rect 79 96 92 99
rect 0 89 107 92
rect 115 87 118 102
rect 0 83 114 86
rect 126 102 152 105
rect 122 80 125 101
rect 135 92 138 95
rect 132 89 138 92
rect 164 93 167 116
rect 164 90 217 93
rect 135 87 138 89
rect 135 84 171 87
rect 203 84 217 87
rect 61 77 200 80
rect 61 31 64 77
rect 91 74 94 77
rect 121 74 124 77
rect 137 74 140 77
rect 167 74 170 77
rect 79 65 82 70
rect 109 65 112 70
rect 73 62 82 65
rect 73 59 76 62
rect 79 59 82 62
rect 103 62 112 65
rect 103 59 106 62
rect 109 59 112 62
rect 149 65 152 70
rect 179 65 182 70
rect 149 62 158 65
rect 149 59 152 62
rect 155 59 158 62
rect 179 62 188 65
rect 179 59 182 62
rect 185 59 188 62
rect 91 52 94 55
rect 121 52 124 55
rect 68 49 129 52
rect 137 52 140 55
rect 167 52 170 55
rect 133 49 193 52
rect 68 41 71 49
rect 80 43 112 46
rect 80 41 83 43
rect 109 41 112 43
rect 121 41 124 49
rect 137 41 140 49
rect 149 43 181 46
rect 149 41 152 43
rect 178 41 181 43
rect 190 41 193 49
rect 95 34 98 36
rect 95 31 141 34
rect 61 28 82 31
rect 79 25 82 28
rect 110 25 113 31
rect 163 27 166 36
rect 197 31 200 77
rect 129 24 166 27
rect 179 28 200 31
rect 68 18 71 21
rect 121 18 124 21
rect 68 15 124 18
rect 129 8 132 24
rect 148 21 151 24
rect 179 21 182 28
rect 137 14 140 17
rect 190 14 193 17
rect 137 11 193 14
rect 203 8 206 84
rect 129 5 206 8
rect 75 0 116 4
<< metal2 >>
rect 71 4 74 129
rect 122 105 125 137
rect 144 86 147 130
rect 130 83 147 86
rect 130 53 133 83
rect 130 4 133 49
rect 120 0 133 4
<< ntransistor >>
rect 27 136 29 139
rect 57 136 59 139
rect 15 118 17 121
rect 27 118 29 121
rect 45 118 47 121
rect 94 123 96 126
rect 104 123 106 126
rect 116 123 118 126
rect 129 123 131 126
rect 136 123 138 126
rect 154 123 156 126
rect 57 118 59 121
rect 86 55 88 58
rect 116 55 118 58
rect 143 55 145 58
rect 173 55 175 58
rect 74 37 76 40
rect 86 37 88 40
rect 104 37 106 40
rect 116 37 118 40
rect 143 37 145 40
rect 155 37 157 40
rect 173 37 175 40
rect 185 37 187 40
<< ptransistor >>
rect 27 150 29 156
rect 57 150 59 156
rect 94 107 96 113
rect 104 107 106 113
rect 116 107 118 113
rect 129 107 131 113
rect 136 107 138 113
rect 154 107 156 113
rect 15 101 17 107
rect 27 101 29 107
rect 45 101 47 107
rect 57 101 59 107
rect 86 69 88 75
rect 116 69 118 75
rect 143 69 145 75
rect 173 69 175 75
rect 74 20 76 26
rect 86 20 88 26
rect 104 20 106 26
rect 116 20 118 26
rect 143 16 145 22
rect 155 16 157 22
rect 173 16 175 22
rect 185 16 187 22
<< polycontact >>
rect 13 136 17 140
rect 43 136 47 140
rect 150 115 154 119
rect 115 102 119 106
rect 92 95 96 99
rect 135 95 139 99
rect 107 89 111 93
rect 128 89 132 93
rect 114 83 118 87
rect 171 83 175 87
rect 72 55 76 59
rect 102 55 106 59
rect 155 55 159 59
rect 185 55 189 59
rect 141 30 145 34
<< ndcontact >>
rect 20 136 24 140
rect 32 136 36 140
rect 50 136 54 140
rect 62 136 66 140
rect 8 118 12 122
rect 20 118 24 122
rect 35 117 39 121
rect 50 118 54 122
rect 88 123 92 127
rect 98 123 102 127
rect 108 123 112 127
rect 122 123 126 127
rect 140 123 144 127
rect 149 123 153 127
rect 157 123 161 127
rect 62 118 66 122
rect 79 55 83 59
rect 91 55 95 59
rect 109 55 113 59
rect 121 55 125 59
rect 136 55 140 59
rect 148 55 152 59
rect 166 55 170 59
rect 178 55 182 59
rect 67 37 71 41
rect 79 37 83 41
rect 94 36 98 40
rect 109 37 113 41
rect 121 37 125 41
rect 136 37 140 41
rect 148 37 152 41
rect 163 36 167 40
rect 178 37 182 41
rect 190 37 194 41
<< pdcontact >>
rect 20 151 24 155
rect 32 151 36 155
rect 50 151 54 155
rect 62 151 66 155
rect 88 108 92 112
rect 98 108 102 112
rect 108 108 112 112
rect 122 108 126 112
rect 140 108 144 112
rect 149 108 153 112
rect 157 108 161 112
rect 8 102 12 106
rect 20 102 24 106
rect 50 102 54 106
rect 62 102 66 106
rect 79 70 83 74
rect 91 70 95 74
rect 109 70 113 74
rect 121 70 125 74
rect 136 70 140 74
rect 148 70 152 74
rect 166 70 170 74
rect 178 70 182 74
rect 67 21 71 25
rect 79 21 83 25
rect 109 21 113 25
rect 121 21 125 25
rect 136 17 140 21
rect 148 17 152 21
rect 178 17 182 21
rect 190 17 194 21
<< m2contact >>
rect 121 137 125 141
rect 70 129 74 133
rect 144 130 148 134
rect 122 101 126 105
rect 129 49 133 53
rect 71 0 75 4
rect 116 0 120 4
<< labels >>
rlabel metal1 213 91 213 91 7 Cout
rlabel metal1 214 85 214 85 7 SUM
rlabel metal1 95 2 95 2 1 gnd
rlabel metal1 81 107 81 107 1 XORB
rlabel metal1 78 138 78 138 1 vdd
rlabel metal1 4 84 4 84 3 A
rlabel metal1 4 91 4 91 3 C
rlabel polysilicon 28 165 28 165 5 B
rlabel polysilicon 58 165 58 165 5 AddSub
<< end >>
