magic
tech scmos
timestamp 1478855084
<< polysilicon >>
rect 3 57 28 60
rect 3 53 6 57
rect 3 46 6 48
rect 3 38 6 42
rect 24 37 28 57
rect 3 24 6 34
rect 3 15 6 19
rect 5 11 6 15
rect 3 6 6 11
rect 3 -2 6 2
<< ndiffusion >>
rect -9 34 -6 38
rect -2 34 3 38
rect 6 34 13 38
rect 17 34 19 38
rect -8 2 -5 6
rect -1 2 3 6
rect 6 2 12 6
rect 16 2 18 6
<< pdiffusion >>
rect -8 49 -6 53
rect -2 49 3 53
rect -8 48 3 49
rect 6 49 13 53
rect 17 49 18 53
rect 6 48 18 49
rect -9 20 -7 24
rect -3 20 3 24
rect -9 19 3 20
rect 6 20 12 24
rect 16 20 17 24
rect 6 19 17 20
<< metal1 >>
rect -6 45 -2 49
rect -16 41 -2 45
rect -6 38 -2 41
rect 3 30 6 64
rect 13 46 17 49
rect 13 42 35 46
rect 13 38 17 42
rect -7 27 6 30
rect -7 24 -3 27
rect 12 16 16 20
rect 24 16 28 32
rect -12 11 1 15
rect 12 12 28 16
rect 12 6 16 12
rect -5 -4 -1 2
<< ntransistor >>
rect 3 34 6 38
rect 3 2 6 6
<< ptransistor >>
rect 3 48 6 53
rect 3 19 6 24
<< polycontact >>
rect 24 32 28 37
rect 1 11 5 15
<< ndcontact >>
rect -6 34 -2 38
rect 13 34 17 38
rect -5 2 -1 6
rect 12 2 16 6
<< pdcontact >>
rect -6 49 -2 53
rect 13 49 17 53
rect -7 20 -3 24
rect 12 20 16 24
<< labels >>
rlabel metal1 -3 -2 -3 -2 1 myGnd
rlabel metal1 -15 43 -15 43 3 myD
rlabel metal1 4 63 4 63 5 myVdd
rlabel metal1 33 43 33 43 7 myQ
rlabel metal1 -9 13 -9 13 1 myC
<< end >>
