* SPICE3 file created from sum.ext - technology: scmos

.option scale=1u

M1000 myVdd myB a_n94_n5# w_n88_66# pfet w=6 l=4
+ ad=378 pd=192 as=42 ps=26 
M1001 myVdd myA a_n59_n5# w_n88_66# pfet w=6 l=4
+ ad=0 pd=0 as=42 ps=26 
M1002 a_32_53# a_n71_30# myVdd w_15_66# pfet w=6 l=4
+ ad=42 pd=26 as=0 ps=0 
M1003 a_64_53# myCin myVdd w_15_66# pfet w=6 l=4
+ ad=42 pd=26 as=0 ps=0 
M1004 myGnd myB a_n94_n5# Gnd nfet w=6 l=4
+ ad=504 pd=264 as=48 ps=28 
M1005 myGnd myA a_n59_n5# Gnd nfet w=6 l=4
+ ad=0 pd=0 as=48 ps=28 
M1006 a_32_53# a_n71_30# myGnd Gnd nfet w=6 l=4
+ ad=48 pd=28 as=0 ps=0 
M1007 a_64_53# myCin myGnd Gnd nfet w=6 l=4
+ ad=48 pd=28 as=0 ps=0 
M1008 a_n90_30# a_n94_n5# myGnd Gnd nfet w=6 l=4
+ ad=162 pd=78 as=0 ps=0 
M1009 a_n71_30# myB a_n90_30# Gnd nfet w=6 l=4
+ ad=72 pd=36 as=0 ps=0 
M1010 a_n90_30# a_n59_n5# a_n71_30# Gnd nfet w=6 l=4
+ ad=0 pd=0 as=0 ps=0 
M1011 myGnd myA a_n90_30# Gnd nfet w=6 l=4
+ ad=0 pd=0 as=0 ps=0 
M1012 a_32_30# a_n71_30# myGnd Gnd nfet w=6 l=4
+ ad=162 pd=78 as=0 ps=0 
M1013 myOut a_32_53# a_32_30# Gnd nfet w=6 l=4
+ ad=72 pd=36 as=0 ps=0 
M1014 a_32_30# myCin myOut Gnd nfet w=6 l=4
+ ad=0 pd=0 as=0 ps=0 
M1015 myGnd a_64_53# a_32_30# Gnd nfet w=6 l=4
+ ad=0 pd=0 as=0 ps=0 
M1016 myVdd a_n94_n5# a_n106_3# w_n109_0# pfet w=7 l=4
+ ad=0 pd=0 as=217 ps=90 
M1017 a_n71_3# myB myVdd w_n109_0# pfet w=7 l=4
+ ad=84 pd=38 as=0 ps=0 
M1018 a_n71_30# a_n59_n5# a_n71_3# w_n109_0# pfet w=7 l=4
+ ad=84 pd=38 as=0 ps=0 
M1019 a_n106_3# myA a_n71_30# w_n109_0# pfet w=7 l=4
+ ad=0 pd=0 as=0 ps=0 
M1020 myOut a_n71_30# a_9_3# w_8_0# pfet w=7 l=4
+ ad=84 pd=38 as=217 ps=90 
M1021 a_48_3# a_32_53# myOut w_8_0# pfet w=7 l=4
+ ad=84 pd=38 as=0 ps=0 
M1022 myVdd myCin a_48_3# w_8_0# pfet w=7 l=4
+ ad=0 pd=0 as=0 ps=0 
M1023 a_9_3# a_64_53# myVdd w_8_0# pfet w=7 l=4
+ ad=0 pd=0 as=0 ps=0 
C0 a_9_3# gnd! 12.0fF
C1 a_n106_3# gnd! 12.0fF
C2 myOut gnd! 14.3fF
C3 a_32_30# gnd! 5.0fF
C4 a_n90_30# gnd! 5.0fF
C5 myGnd gnd! 48.3fF
C6 a_64_53# gnd! 20.8fF
C7 a_32_53# gnd! 19.7fF
C8 a_n59_n5# gnd! 19.7fF
C9 myVdd gnd! 87.2fF
C10 a_n94_n5# gnd! 20.8fF
C11 myCin gnd! 20.9fF
C12 a_n71_30# gnd! 41.0fF
C13 myA gnd! 20.9fF
C14 myB gnd! 20.9fF


.include ../usc-spice.usc-spice

Vgnd1 myGnd 0 DC 0V
Vgnd2 gnd! 0 DC 0V

VVdd myVdd 0 DC 2.8V

Vin1 myA 0 pulse(0 2.8v 0ns 0.1ns 0.1ns 64ns 128ns)
Vin2 myB 0 pulse(0 2.8v 0ns 0.1ns 0.1ns 128ns 256ns)
Vin3 myCin 0 pulse(0 2.8v 0ns 0.1ns 0.1ns 256ns 512ns)

.tran 1ns 1000ns
.probe
.control
run
plot myA myB+4 myCin+8 myOut+12
.endc
.end
