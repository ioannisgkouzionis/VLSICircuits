magic
tech scmos
timestamp 1478776710
<< polysilicon >>
rect -2 17 1 19
rect 10 17 13 19
rect 31 17 34 19
rect -2 -26 1 10
rect 10 -26 13 10
rect 31 -7 34 10
rect 32 -13 34 -7
rect 31 -26 34 -13
rect -2 -36 1 -32
rect 10 -36 13 -32
rect 31 -36 34 -32
<< ndiffusion >>
rect -12 -27 -2 -26
rect -12 -31 -9 -27
rect -5 -31 -2 -27
rect -12 -32 -2 -31
rect 1 -32 10 -26
rect 13 -27 20 -26
rect 13 -31 15 -27
rect 19 -31 20 -27
rect 13 -32 20 -31
rect 23 -27 31 -26
rect 23 -31 25 -27
rect 29 -31 31 -27
rect 23 -32 31 -31
rect 34 -27 46 -26
rect 34 -31 40 -27
rect 44 -31 46 -27
rect 34 -32 46 -31
<< pdiffusion >>
rect -8 15 -2 17
rect -8 11 -7 15
rect -3 11 -2 15
rect -8 10 -2 11
rect 1 15 10 17
rect 1 11 4 15
rect 8 11 10 15
rect 1 10 10 11
rect 13 15 31 17
rect 13 11 19 15
rect 23 11 31 15
rect 13 10 31 11
rect 34 15 43 17
rect 34 11 36 15
rect 40 11 43 15
rect 34 10 43 11
<< metal1 >>
rect -7 20 23 23
rect -7 15 -3 20
rect 19 15 23 20
rect 4 3 8 11
rect 36 8 40 11
rect 36 5 51 8
rect -15 -4 -7 2
rect 4 -1 19 3
rect 15 -7 19 -1
rect -15 -13 5 -7
rect 15 -13 27 -7
rect 15 -27 19 -13
rect 40 -27 44 5
rect -9 -41 -5 -31
rect 25 -41 29 -31
rect -9 -44 29 -41
rect -9 -47 -5 -44
<< ntransistor >>
rect -2 -32 1 -26
rect 10 -32 13 -26
rect 31 -32 34 -26
<< ptransistor >>
rect -2 10 1 17
rect 10 10 13 17
rect 31 10 34 17
<< polycontact >>
rect -7 -4 -2 2
rect 5 -13 10 -7
rect 27 -13 32 -7
<< ndcontact >>
rect -9 -31 -5 -27
rect 15 -31 19 -27
rect 25 -31 29 -27
rect 40 -31 44 -27
<< pdcontact >>
rect -7 11 -3 15
rect 4 11 8 15
rect 19 11 23 15
rect 36 11 40 15
<< labels >>
rlabel metal1 -13 -1 -13 -1 3 myB
rlabel metal1 -12 -10 -12 -10 3 myA
rlabel metal1 -5 21 -5 21 5 myVdd
rlabel metal1 49 7 49 7 7 myOut
rlabel metal1 -7 -46 -7 -46 1 myGnd
<< end >>
