* SPICE3 file created from and.ext - technology: scmos

.option scale=1u

M1000 a_1_10# myB myVdd Vdd pfet w=7 l=3
+ ad=63 pd=32 as=168 ps=76 
M1001 myVdd myA a_1_10# Vdd pfet w=7 l=3
+ ad=0 pd=0 as=0 ps=0 
M1002 myOut a_1_10# myVdd Vdd pfet w=7 l=3
+ ad=63 pd=32 as=0 ps=0 
M1003 a_1_n32# myB myGnd Gnd nfet w=6 l=3
+ ad=54 pd=30 as=108 ps=60 
M1004 a_1_10# myA a_1_n32# Gnd nfet w=6 l=3
+ ad=42 pd=26 as=0 ps=0 
M1005 myOut a_1_10# myGnd Gnd nfet w=6 l=3
+ ad=72 pd=36 as=0 ps=0 
C0 myGnd gnd! 9.3fF
C1 myOut gnd! 8.3fF
C2 myVdd gnd! 5.4fF
C3 a_1_10# gnd! 25.2fF
C4 myA gnd! 19.8fF
C5 myB gnd! 17.3fF

.include ../usc-spice.usc-spice

Vgnd1 myGnd 0 DC 0V
Vgnd2 gnd! 0 DC 0V

VVdd myVdd 0 DC 2.8V

Vin1 myA 0 pulse(0 2.8v 0ns 0.1ns 0.1ns 64ns 128ns)
Vin2 myB 0 pulse(0 2.8v 0ns 0.1ns 0.1ns 128ns 256ns)

.tran 1ns 1000ns
.probe
.control
run
plot myA myB+4 myOut+8
.endc
.end