magic
tech scmos
timestamp 1480950362
<< polysilicon >>
rect 4 13 6 15
<< metal1 >>
rect 0 29 40 32
rect 0 23 3 29
rect 37 23 40 29
rect 11 13 39 16
rect 48 14 62 17
rect 0 3 3 7
rect 37 3 40 8
rect 0 0 40 3
<< polycontact >>
rect 39 13 43 17
use inverter  inverter_0
timestamp 1351319193
transform 1 0 5 0 1 13
box -5 -10 7 15
use inverter  inverter_1
timestamp 1351319193
transform 1 0 42 0 1 13
box -5 -10 7 15
<< labels >>
rlabel metal1 20 31 20 31 5 Vdd!
rlabel metal1 20 1 20 1 1 GND!
rlabel polysilicon 5 14 5 14 3 Vin
rlabel metal1 13 15 13 15 1 Vout
rlabel metal1 61 15 61 15 7 out
<< end >>
